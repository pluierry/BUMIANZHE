`define Temp_BJ 40'h781c0712a0 //����
`define Temp_TJ 40'h7beef752e0 //���
`define Temp_HB 40'h7edce779f1 //�ӱ�
`define Temp_SX 40'hfbfee53a42 //ɽ��
`define Temp_NM 40'hfffffff7a5 //����
`define Temp_LN 40'h7844211387 //����
`define Temp_JL 40'h3fc84743c0 //����
`define Temp_HL 40'h7bdec77fa1 //������
`define Temp_SH 40'h7be254e300 //�Ϻ�
`define Temp_JS 40'h7b98eded44 //����
`define Temp_ZZ 40'hfb28f77b8c //�㽭
`define Temp_AH 40'h7f7f8ffae1 //����
`define Temp_FJ 40'h7d7fffde62 //����
`define Temp_JX 40'h7fbfefffe5 //����
`define Temp_SD 40'h7f9ee7b9c2 //ɽ��
`define Temp_NH 40'h7bdff7b9e0 //����
`define Temp_UB 40'hffdebfacc8 //����
`define Temp_UN 40'hfb6ed7f6e1 //����
`define Temp_GD 40'h7bdfffb846 //�㶫 
`define Temp_GX 40'h7fc5ff09c0 //����
`define Temp_HN 40'h7a0fd3b964 //����
`define Temp_CC 40'h7bbaf7ffa6 //����
`define Temp_SC 40'h7b5ad296a0 //�Ĵ�
`define Temp_GZ 40'hffff87e7c2 //����
`define Temp_YN 40'hf9aef7fec1 //����
`define Temp_XZ 40'h7bfdfffbe5 //����
`define Temp_AX 40'hffffeffa81 //����
`define Temp_GS 40'h7fc4a509c0 //����
`define Temp_QS 40'h7bbee77a42 //�ຣ
`define Temp_NX 40'h3fc3f21088 //����
`define Temp_XJ 40'h7b38f77b80 //�½�

 
`define A     "A"
`define B     "B"
`define C     "C"
`define D     "D"
`define E     "E"
`define F     "F"
`define G     "G"
`define H     "H"
`define I     "I"
`define J     "J"
`define K     "K"
`define L     "L"
`define M     "M"
`define N     "N"
`define P     "P"
`define Q     "Q"
`define R     "R"
`define S     "S"
`define T     "T"
`define U     "U"
`define V     "V"
`define W     "W"
`define X     "X"
`define Y     "Y"
`define Z     "Z"
