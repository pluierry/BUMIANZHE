`define Temp_A 40'h3b1ce57bf1
`define Temp_B 40'hfcf7e9cf7c
`define Temp_C 40'h7e6108432e
`define Temp_D 40'hfce318c63f
`define Temp_E 40'hfc21ec421f
`define Temp_F 40'hfe21ec4210
`define Temp_G 40'h7c6179c62e
`define Temp_H 40'hfc63bdc631
`define Temp_I 40'hf98c6310df
`define Temp_J 40'h084210876e
`define Temp_K 40'hfcbded4e71
`define Temp_L 40'hfe318c631f
`define Temp_M 40'hfffff8c631
`define Temp_N 40'hfe7bfbee7b
`define Temp_P 40'hfef3fe6318
`define Temp_Q 40'h7c6318c7ef
`define Temp_R 40'hfc63bf5a53
`define Temp_S 40'h7ee0e1876e
`define Temp_T 40'hf908421084
`define Temp_U 40'h746318c631
`define Temp_V 40'hfef4a73984
`define Temp_W 40'h5295ffd6b1
`define Temp_X 40'hfa9c423953
`define Temp_Y 40'hfa9c423184
`define Temp_Z 40'h78c462231f

`define Temp_0 40'h7ee318c76e
`define Temp_1 40'hffffffffff
`define Temp_2 40'h7cc622331f
`define Temp_3 40'hf888e1876e
`define Temp_4 40'h198ca56fe2
`define Temp_5 40'hfe31e1876e
`define Temp_6 40'h3911cfc72e
`define Temp_7 40'hf8c4231084
`define Temp_8 40'h7e72edc76e
`define Temp_9 40'h7ee3f3988c 
 
`define A     "A"
`define B     "B"
`define C     "C"
`define D     "D"
`define E     "E"
`define F     "F"
`define G     "G"
`define H     "H"
`define I     "I"
`define J     "J"
`define K     "K"
`define L     "L"
`define M     "M"
`define N     "N"
`define P     "P"
`define Q     "Q"
`define R     "R"
`define S     "S"
`define T     "T"
`define U     "U"
`define V     "V"
`define W     "W"
`define X     "X"
`define Y     "Y"
`define Z     "Z"

`define NUM0 "0"
`define NUM1 "1"
`define NUM2 "2"
`define NUM3 "3"
`define NUM4 "4"
`define NUM5 "5"
`define NUM6 "6"
`define NUM7 "7"
`define NUM8 "8"
`define NUM9 "9"
